--Nama      : Rifki Afriadi
--NIM       : 13223049
--Rombongan : C
--Kelompok  : 7
--Percobaan : 2B
--Tanggal   : 14/10/2024


--Deskripsi
--Fungsi : Mengubah bilangan BCD satu digit(4bit) menjadi bentuk seven segment satu digit
--Input : SW (4 digit)
--Output : HEX1(4 BIT)

LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.numeric_std.all;
ENTITY bcd IS PORT (
 SW : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
 HEX1 : OUT STD_LOGIC_VECTOR (1 TO 7));
END bcd;
ARCHITECTURE behavioral OF bcd IS
CONSTANT NOL : STD_LOGIC_VECTOR(3 DOWNTO 0) := "0000";
CONSTANT SATU : STD_LOGIC_VECTOR(3 DOWNTO 0) := "0001";
CONSTANT DUA : STD_LOGIC_VECTOR(3 DOWNTO 0) := "0010";
CONSTANT TIGA : STD_LOGIC_VECTOR(3 DOWNTO 0) := "0011";
CONSTANT EMPAT : STD_LOGIC_VECTOR(3 DOWNTO 0) := "0100";
CONSTANT LIMA : STD_LOGIC_VECTOR(3 DOWNTO 0) := "0101";
CONSTANT ENAM : STD_LOGIC_VECTOR(3 DOWNTO 0) := "0110";
CONSTANT TUJUH : STD_LOGIC_VECTOR(3 DOWNTO 0) := "0111";
CONSTANT DELAPAN : STD_LOGIC_VECTOR(3 DOWNTO 0) := "1000";
CONSTANT SEMBILAN: STD_LOGIC_VECTOR(3 DOWNTO 0) := "1001";
BEGIN
PROCESS(SW)
BEGIN
CASE SW IS
WHEN NOL => HEX1 <= NOT "1111110";
WHEN SATU => HEX1 <= NOT "0110000";
WHEN DUA => HEX1 <= NOT "1101101";
WHEN TIGA => HEX1 <= NOT "1111001";
WHEN EMPAT => HEX1 <= NOT "0110011";
WHEN LIMA => HEX1 <= NOT "1011011";
WHEN ENAM => HEX1 <= NOT "1011111";
WHEN TUJUH => HEX1 <= NOT "1110000";
WHEN DELAPAN => HEX1 <= NOT "1111111";
WHEN SEMBILAN => HEX1 <= NOT "1110011";
WHEN OTHERS => HEX1 <=  "0000000";
END CASE;
END PROCESS;
END behavioral;